// Global include file for register interface and AXI typedef structures
// Created for particular use in development process
//

`include "register_interface/typedef.svh"
`include "axi/typedef.svh"
`include "axi_pkg.sv"

`ifndef GLOBAL_TYPEDEF_SVH
`define GLOBAL_TYPEDEF_SVH

typedef logic [64-1:0]  addr_t;
typedef logic [64-1:0]  data_t;
typedef logic [8-1:0]   strb_t;

// Define reg_req_t and reg_rsp_t structs
`REG_BUS_TYPEDEF_ALL(iommu_reg, addr_t, data_t, strb_t)

`endif
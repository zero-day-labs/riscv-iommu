// Copyright © 2024 Manuel Rodríguez & Zero-Day Labs, Lda.
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1

// Licensed under the Solderpad Hardware License v 2.1 (the “License”); 
// you may not use this file except in compliance with the License, 
// or, at your option, the Apache License version 2.0. 
// You may obtain a copy of the License at https://solderpad.org/licenses/SHL-2.1/.
// Unless required by applicable law or agreed to in writing, 
// any work distributed under the License is distributed on an “AS IS” BASIS, 
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
// See the License for the specific language governing permissions and limitations under the License.
//
// Author: Manuel Rodríguez <manuel.cederog@gmail.com>
// Date: 21/05/2024
// Acknowledges: SSRC - Technology Innovation Institute (TII)
//
// Description: Slave module to ignore requests within the IOMMU and provide completions.

module rv_iommu_ign_slv #(
    /// AXI ID Width
    parameter int unsigned          AxiIdWidth  = 0,
    /// Response generated by the slave
    parameter axi_pkg::resp_t       Resp        = axi_pkg::RESP_OKAY,
    /// Data response width, gets zero extended or truncated to r.data
    parameter int unsigned          RespWidth   = 32'd64,
    /// Hexvalue for data return value
    parameter logic [RespWidth-1:0] RespData    = 64'h0,
    /// AXI Full request struct type
    parameter type                  axi_req_t   = logic,
    /// AXI Full response struct type
    parameter type                  axi_rsp_t   = logic
) (
    input  logic        clk_i,
    input  logic        rst_ni,
    
    input  axi_req_t    ignore_req_i,
    output axi_rsp_t    ignore_resp_o
);

    logic [(AxiIdWidth-1):0]    b_id_q, b_id_n;
    logic [(AxiIdWidth-1):0]    r_id_q, r_id_n;
    logic [7:0]                 r_counter_q, r_counter_n;

    logic   ign_aw_ready_q, ign_aw_ready_n;
    logic   ign_w_ready_q,  ign_w_ready_n;
    logic   ign_b_valid_q,  ign_b_valid_n;
    logic   ign_ar_ready_q, ign_ar_ready_n;
    logic   ign_r_valid_q,  ign_r_valid_n;

    always_comb begin : ignore_req_comb

        // Set output signals
        ignore_resp_o.aw_ready  = ign_aw_ready_q;
        ignore_resp_o.w_ready   = ign_w_ready_q;
        ignore_resp_o.b_valid   = ign_b_valid_q;
        ignore_resp_o.ar_ready  = ign_ar_ready_q;
        ignore_resp_o.r_valid   = ign_r_valid_q;

        ignore_resp_o.b.id      = b_id_q;
        ignore_resp_o.b.resp    = Resp;
        ignore_resp_o.b.user    = '0;

        ignore_resp_o.r.id      = r_id_q;
        ignore_resp_o.r.data    = RespData;
        ignore_resp_o.r.resp    = Resp;
        ignore_resp_o.r.last    = (r_counter_q == '0) & ign_r_valid_q;
        ignore_resp_o.r.user    = '0;

        // Default assignments
        b_id_n          = b_id_q;
        r_id_n          = r_id_q;
        r_counter_n     = r_counter_q;

        ign_aw_ready_n  = 1'b0;
        ign_w_ready_n   = ign_w_ready_q;
        ign_b_valid_n   = ign_b_valid_q;
        ign_ar_ready_n  = 1'b0;
        ign_r_valid_n   = ign_r_valid_q;

        // Read transaction
        if (ignore_req_i.ar_valid) begin
            
            // Save ARID
            r_id_n          = ignore_req_i.ar.id;
            // Save number of read transfers
            r_counter_n     = ignore_req_i.ar.len;

            if (!ign_ar_ready_q)
                // Set ARREADY
                ign_ar_ready_n  = 1'b1;
            else
                // Set RVALID when ARREADY is set by IOMMU
                ign_r_valid_n = 1'b1;
        end

        // Send requested beats
        if (ign_r_valid_q && ignore_req_i.r_ready) begin
            
            // Clear RVALID when counter reaches zero    
            if (r_counter_q == '0)
                ign_r_valid_n = 1'b0;
            else
                // Decrement counter
                r_counter_n  = r_counter_q - 1;
        end

        // Write transaction
        if (ignore_req_i.aw_valid) begin
            // Set AWREADY
            if (!ign_aw_ready_q)
                ign_aw_ready_n  = 1'b1;
            // Save AWID
            b_id_n          = ignore_req_i.aw.id;
        end

        // Receive all write beats
        if (ignore_req_i.w_valid) begin
            // Set WREADY after WVALID is set by master
            ign_w_ready_n = 1'b1;

            if (ignore_req_i.w.last && ign_w_ready_q) begin
                // Clear WREADY when WLAST is set by master
                ign_w_ready_n = 1'b0;
                // Set BVALID
                ign_b_valid_n = 1'b1;
            end
        end 
        
        // Clear BVALID when master sets BREADY
        if (ign_b_valid_q && ignore_req_i.b_ready)
            ign_b_valid_n = 1'b0;

    end : ignore_req_comb

    always_ff @( posedge clk_i or negedge rst_ni ) begin : ignore_req_ff

        if (~rst_ni) begin
            b_id_q          <= '0;
            r_id_q          <= '0;
            r_counter_q     <= '0;

            ign_aw_ready_q  <= 1'b0;
            ign_w_ready_q   <= 1'b0;
            ign_b_valid_q   <= 1'b0;
            ign_ar_ready_q  <= 1'b0;
            ign_r_valid_q   <= 1'b0;
        end

        else begin
            b_id_q          <= b_id_n;
            r_id_q          <= r_id_n;
            r_counter_q     <= r_counter_n;
            
            ign_aw_ready_q  <= ign_aw_ready_n;
            ign_w_ready_q   <= ign_w_ready_n;
            ign_b_valid_q   <= ign_b_valid_n;
            ign_ar_ready_q  <= ign_ar_ready_n;
            ign_r_valid_q   <= ign_r_valid_n;
        end
    end : ignore_req_ff
endmodule
// Copyright © 2023 Manuel Rodríguez & Zero-Day Labs, Lda.
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1

// Licensed under the Solderpad Hardware License v 2.1 (the “License”); 
// you may not use this file except in compliance with the License, 
// or, at your option, the Apache License version 2.0. 
// You may obtain a copy of the License at https://solderpad.org/licenses/SHL-2.1/.
// Unless required by applicable law or agreed to in writing, 
// any work distributed under the License is distributed on an “AS IS” BASIS, 
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
// See the License for the specific language governing permissions and limitations under the License.
//
// Author: Manuel Rodríguez <manuel.cederog@gmail.com>
// Date: 06/02/2023
// Acknowledges: SSRC - Technology Innovation Institute (TII)
//
// Description: RISC-V IOMMU Translation Logic Wrapper.
//              Encompasses all modules involved in the address translation 
//              process and report of translation faults.
//              Process Context support: NO
//              MSI Translation support: YES

//! NOTES:
/*
    - For now, req_trans_i must be hold high for the entire translation process (whenever walks are needed). If it is cleared, 
      IOTLB hit signal is also cleared even if it has a valid translation. Further on, input signals may be propagated to achieve 
      a stronger implementation (+ HW cost).
*/

module rv_iommu_tw_sv39x4_msi #(

    parameter int unsigned  IOTLB_ENTRIES       = 4,
    parameter int unsigned  DDTC_ENTRIES        = 4,

    /// AXI Full request struct type
    parameter type  axi_req_t       = logic,
    /// AXI Full response struct type
    parameter type  axi_rsp_t       = logic
) (
    input  logic    clk_i,
    input  logic    rst_ni,

    // Trigger translation
    input  logic    req_trans_i,

    // Translation request data
    input  logic [23:0]                     did_i,      // device_id associated with the transaction
    input  logic [riscv::VLEN-1:0]          iova_i,     // IOVA
    output logic [15:0]                     gscid_o,    // GSCID
    output logic [19:0]                     pscid_o,    // PSCID
    
    input  logic [rv_iommu::TTYP_LEN-1:0]   trans_type_i,   // transaction type

    // AXI ports directed to Data Structures Interface
    // CDW
    input  axi_rsp_t   cdw_axi_resp_i,
    output axi_req_t    cdw_axi_req_o,
    // PTW
    input  axi_rsp_t   ptw_axi_resp_i,
    output axi_req_t    ptw_axi_req_o,

    // From Regmap
    input  rv_iommu_reg_pkg::iommu_reg2hw_capabilities_reg_t   capabilities_i,
    input  rv_iommu_reg_pkg::iommu_reg2hw_fctl_reg_t           fctl_i,
    input  rv_iommu_reg_pkg::iommu_reg2hw_ddtp_reg_t           ddtp_i,

    // Request status and output data
    output logic                        trans_valid_o,      // Translation completed
    output logic [riscv::PLEN-1:0]      spaddr_o,           // Translated address
    output logic                        is_msi_o,           // Indicate whether the translated address is an MSI address
    // Error
    output logic                                trans_error_o,      // Translation error
    output logic                                report_fault_o,     // The fault must be reported through the FQ
    output logic [(rv_iommu::CAUSE_LEN-1):0]    cause_code_o,       // Fault code defined by translation logic
    output logic                                is_guest_pf_o,      // a guest page fault occurred in the PTW
    output logic                                is_implicit_o,      // Guest page fault caused by implicit access for 1st-stage addr translation
    output logic [riscv::SVX-1:0]               bad_gpaddr_o,       // to report bits [63:2] of the GPA in case of a Guest Page Fault
    input  logic                                msi_write_error_i,  // An error occurred when writing an MSI generated by the IOMMU

    // to HPM
    output logic                        iotlb_miss_o,       // IOTLB miss happened
    output logic                        ddt_walk_o,         // DDT walk triggered
    output logic                        pdt_walk_o,         // PDT walk triggered
    output logic                        s1_ptw_o,           // first-stage PT walk triggered
    output logic                        s2_ptw_o,           // second-stage PT walk triggered

    // IOATC Invalidation control (from CQ Handler to IOATC)
    // DDTC Invalidation
    input  logic                        flush_ddtc_i,   // Flush DDTC
    input  logic                        flush_dv_i,     // Indicates if device_id is valid
    input  logic [23:0]                 flush_did_i,    // device_id to tag entries to be flushed
    // IOTLB Invalidation
    input  logic                        flush_vma_i,    // Flush first-stage PTEs cached entries in IOTLB
    input  logic                        flush_gvma_i,   // Flush second-stage PTEs cached entries in IOTLB 
    input  logic                        flush_av_i,     // Address valid
    input  logic                        flush_gv_i,     // GSCID valid
    input  logic                        flush_pscv_i,   // PSCID valid
    input  logic [riscv::GPPNW-1:0]     flush_vpn_i,    // IOVA to tag entries to be flushed
    input  logic [15:0]                 flush_gscid_i,  // GSCID (Guest physical address space identifier) to tag entries to be flushed
    input  logic [19:0]                 flush_pscid_i   // PSCID (Guest virtual address space identifier) to tag entries to be flushed
);

    // DDTC
    logic                       ddtc_access;
    rv_iommu::dc_ext_t          ddtc_lu_content;
    logic                       ddtc_lu_hit;

    // IOTLB
    logic                       iotlb_access;
    logic [riscv::GPLEN-1:0]    iotlb_lu_gpaddr;
    riscv::pte_t                iotlb_lu_1S_content;
    riscv::pte_t                iotlb_lu_2S_content;
    logic                       iotlb_lu_1S_2M;
    logic                       iotlb_lu_1S_1G;
    logic                       iotlb_lu_2S_2M;
    logic                       iotlb_lu_2S_1G;
    logic                       iotlb_lu_is_msi;
    logic                       iotlb_lu_hit;

    // Bare translation signaled by PTW
    logic is_bare_translation;

    // PTW error
    logic ptw_error;
    logic [(rv_iommu::CAUSE_LEN-1):0]  ptw_cause_code;

    // CDW error
    logic cdw_error;
    logic [(rv_iommu::CAUSE_LEN-1):0]  cdw_cause_code;

    // Address translation parameters
    logic en_1S, en_2S;
    logic [15:0] gscid;
    logic [19:0] pscid;
    logic [riscv::PPNW-1:0] iohgatp_ppn, iosatp_ppn;

    // To check whether first and second-stage translation modes are Bare
    logic first_stage_is_bare, second_stage_is_bare;
    assign first_stage_is_bare  =   (ddtc_lu_content.fsc.mode == 4'b0000);
    assign second_stage_is_bare =   (ddtc_lu_content.iohgatp.mode == 4'b0000);

    // To determine if current DC enables MSI translation
    logic msi_enabled;
    assign msi_enabled = (ddtc_lu_content.msiptp.mode != 4'b0000);

    // To determine if request is translated or untranslated
    logic is_translated;
    assign is_translated = (!trans_type_i[3] && trans_type_i[2]);

    // To determine if request is a PCIe ATS TR
    logic is_pcie_tr_req;
    assign is_pcie_tr_req = (trans_type_i == rv_iommu::PCIE_ATS_TRANS_REQ);

    // To determine if transaction is a store
    logic is_store;
    assign is_store = ((&trans_type_i[1:0] == 1'b1) && (!trans_type_i[3]));

    // To determine if transaction is read-for-execute
    logic is_rx;
    assign is_rx = (!trans_type_i[3] && !trans_type_i[1] && trans_type_i[0]);

    // Efective iohgatp.ppn field to introduce in the PTW. May need to be forwarded by the CDW
    logic [riscv::PPNW-1:0] ptw_iohgatp_ppn;
    assign ptw_iohgatp_ppn = iohgatp_ppn;

    // To select en_1S and en_2S source
    logic   ptw_en_1S, ptw_en_2S;
    assign  ptw_en_1S = en_1S;
    assign  ptw_en_2S = en_2S;

    // Set for faults occurred before DDTC lookup
    logic   report_always;

    // Error/fault signaling according to the spec
    logic   trans_error;
    assign  trans_error_o = trans_error;  // The requesting device needs to know if an error occurred

    logic [(rv_iommu::CAUSE_LEN-1):0]  cause_code;  // Fault code as defined by IOMMU and Priv Spec
    assign cause_code_o = cause_code;

    // To indicate whether the occurring fault has to be reported according to DC.tc.DTF and the fault source
    // If DC.tc.DTF=1, only faults occurred before finding the corresponding DC should be reported
    assign  report_fault_o    = (((ddtc_lu_hit & !ddtc_lu_content.tc.dtf) | 
                                  (report_always | msi_write_error_i | cdw_error)) & trans_error);
                                  
    // Guest page fault occurred during implicit 2nd-stage translation for 1st-stage translation
    logic   ptw_error_2S_int;
    assign  is_implicit_o = (ptw_error_2S_int);

    // HPM event indicators
    logic cdw_active, ptw_active;
    assign iotlb_miss_o = iotlb_access & (~iotlb_lu_hit);
    assign ddt_walk_o   = cdw_active;
    assign pdt_walk_o   = 1'b0;
    assign s1_ptw_o     = ptw_active & (ptw_en_1S);
    assign s2_ptw_o     = ptw_active & (ptw_en_2S);
    assign gscid_o      = gscid;
    assign pscid_o      = pscid;


    // Update wires
    logic                       ddtc_update;
    logic [23:0]                ddtc_up_did;
    rv_iommu::dc_ext_t          ddtc_up_content;

    logic                       iotlb_update;
    logic                       iotlb_up_1S_2M;
    logic                       iotlb_up_1S_1G;
    logic                       iotlb_up_2S_2M;
    logic                       iotlb_up_2S_1G;
    logic                       iotlb_up_is_msi;
    logic [riscv::GPPNW-1:0]    iotlb_up_vpn;
    logic [19:0]                iotlb_up_pscid;
    logic [15:0]                iotlb_up_gscid;
    riscv::pte_t                iotlb_up_1S_content;
    riscv::pte_t                iotlb_up_2S_content;

    //# Device Directory Table Cache
    rv_iommu_ddtc #(
        .DDTC_ENTRIES       (DDTC_ENTRIES),
        .dc_t               (rv_iommu::dc_ext_t)
    ) i_rv_iommu_ddtc (
        .clk_i              (clk_i          ),  // Clock
        .rst_ni             (rst_ni         ),  // Asynchronous reset active low

        .flush_i            (flush_ddtc_i   ),  // IODIR.INVAL_DDT
        .flush_dv_i         (flush_dv_i     ),  // device_id valid
        .flush_did_i        (flush_did_i    ),  // device_id to be flushed

        // Update signals
        .update_i           (ddtc_update    ),  // update flag
        .up_did_i           (ddtc_up_did    ),  // device ID to be updated
        .up_content_i       (ddtc_up_content),  // DC to be inserted

        // Lookup signals
        .lookup_i           (ddtc_access    ),  // lookup flag
        .lu_did_i           (did_i          ),  // device_id to look for 
        .lu_content_o       (ddtc_lu_content),  // DC found in DDTC
        .lu_hit_o           (ddtc_lu_hit    )   // hit flag
    );

    //# IOTLB: Address Translation Cache
    rv_iommu_iotlb_sv39x4_msi #(
        .IOTLB_ENTRIES      (IOTLB_ENTRIES)
    ) i_rv_iommu_iotlb_sv39x4_msi (
        .clk_i              (clk_i      ),  // Clock
        .rst_ni             (rst_ni     ),  // Asynchronous reset active low

        // Flush signals
        .flush_vma_i        (flush_vma_i        ),  // IOTINVAL.VMA
        .flush_gvma_i       (flush_gvma_i       ),  // IOTINVAL.GVMA
        .flush_av_i         (flush_av_i         ),  // ADDR valid
        .flush_gv_i         (flush_gv_i         ),  // GSCID valid
        .flush_pscv_i       (flush_pscv_i       ),  // PSCID valid
        .flush_vpn_i        (flush_vpn_i        ),  // VPN to be flushed
        .flush_gscid_i      (flush_gscid_i      ),  // GSCID identifier to be flushed (VM identifier)
        .flush_pscid_i      (flush_pscid_i      ),  // PSCID identifier to be flushed (address space identifier)

        // Update signals
        .update_i           (iotlb_update       ),
        .up_1S_2M_i         (iotlb_up_1S_2M     ),
        .up_1S_1G_i         (iotlb_up_1S_1G     ),
        .up_2S_2M_i         (iotlb_up_2S_2M     ),
        .up_2S_1G_i         (iotlb_up_2S_1G     ),
        .up_is_msi_i        (iotlb_up_is_msi    ),
        .up_vpn_i           (iotlb_up_vpn       ),
        .up_pscid_i         (iotlb_up_pscid     ),
        .up_gscid_i         (iotlb_up_gscid     ),
        .up_1S_content_i    (iotlb_up_1S_content),
        .up_2S_content_i    (iotlb_up_2S_content),

        // Lookup signals
        .lookup_i           (iotlb_access       ),  // lookup flag
        .lu_iova_i          (iova_i             ),  // IOVA to look for 
        .lu_pscid_i         (pscid              ),  // PSCID to look for
        .lu_gscid_i         (gscid              ),  // GSCID to look for
        .lu_gpaddr_o        (iotlb_lu_gpaddr    ),  // GPA to return in case of an exception
        .lu_1S_content_o    (iotlb_lu_1S_content),  // first-stage PTE (GPA PPN)
        .lu_2S_content_o    (iotlb_lu_2S_content),  // second-stage PTE (SPA PPN)
        .lu_1S_2M_o         (iotlb_lu_1S_2M     ),
        .lu_1S_1G_o         (iotlb_lu_1S_1G     ),
        .lu_2S_2M_o         (iotlb_lu_2S_2M     ),
        .lu_2S_1G_o         (iotlb_lu_2S_1G     ),
        .lu_is_msi_o        (iotlb_lu_is_msi    ),  // IOTLB entry contains a GPA associated with a guest vIMSIC
        .en_1S_i            (en_1S              ),  // first-stage enabled
        .en_2S_i            (en_2S              ),  // second-stage enabled
        .lu_hit_o           (iotlb_lu_hit       )   // hit flag
    );

    //# Page Table Walker
    rv_iommu_ptw_sv39x4_msi #(
        .axi_req_t          (axi_req_t ),
        .axi_rsp_t          (axi_rsp_t )
    ) i_rv_iommu_ptw_sv39x4_msi (
        .clk_i                  (clk_i              ),  // Clock
        .rst_ni                 (rst_ni             ),  // Asynchronous reset active low
        
        // Error signaling
        .ptw_active_o           (ptw_active         ),  // Set when PTW is walking memory
        .ptw_error_o            (ptw_error          ),  // set when an error occurred (excluding access errors)
        .ptw_error_2S_o         (is_guest_pf_o      ),  // set when the fault occurred in stage 2
        .ptw_error_2S_int_o     (ptw_error_2S_int   ),  // set when fault occurred during an implicit access for 1st-stage translation
        .cause_code_o           (ptw_cause_code     ),

        .en_1S_i                (ptw_en_1S          ),  // Enable signal for stage 1 translation. Defined by DC/PC
        .en_2S_i                (ptw_en_2S          ),  // Enable signal for stage 2 translation. Defined by DC only
        .is_store_i             (is_store           ),  // Indicate whether this translation was triggered by a store or a load
        .is_rx_i                (is_rx              ),  // Read-for-execute

        // PTW AXI Master memory interface
        .mem_resp_i             (ptw_axi_resp_i     ),  // Response port from memory
        .mem_req_o              (ptw_axi_req_o      ),  // Request port to memory

        // to IOTLB, update logic
        .update_o               (iotlb_update       ),
        .up_1S_2M_o             (iotlb_up_1S_2M     ),
        .up_1S_1G_o             (iotlb_up_1S_1G     ),
        .up_2S_2M_o             (iotlb_up_2S_2M     ),
        .up_2S_1G_o             (iotlb_up_2S_1G     ),
        .up_is_msi_o            (iotlb_up_is_msi    ),
        .up_vpn_o               (iotlb_up_vpn       ),
        .up_pscid_o             (iotlb_up_pscid     ),
        .up_gscid_o             (iotlb_up_gscid     ),
        .up_1S_content_o        (iotlb_up_1S_content),
        .up_2S_content_o        (iotlb_up_2S_content),

        // IOTLB tags
        .req_iova_i             (iova_i             ),
        .pscid_i                (pscid              ),
        .gscid_i                (gscid              ),

        // MSI translation
        .msi_en_i               (msi_enabled                                ),
        .msiptp_ppn_i           (ddtc_lu_content.msiptp.ppn                 ),
        .msi_addr_mask_i        (ddtc_lu_content.msi_addr_mask.mask         ),
        .msi_addr_pattern_i     (ddtc_lu_content.msi_addr_pattern.pattern   ),
        .bare_translation_o     (is_bare_translation                        ),     // both stages are in bare mode and address is not MSI

        // from IOTLB, to monitor misses
        .iotlb_access_i         (iotlb_access       ),
        .iotlb_hit_i            (iotlb_lu_hit       ),

        // from DC/PC
        .iosatp_ppn_i           (iosatp_ppn         ),  // ppn from iosatp
        .iohgatp_ppn_i          (ptw_iohgatp_ppn    ),  // ppn from iohgatp (may be forwarded by the CDW)

        .bad_gpaddr_o           (bad_gpaddr_o       )   // to return the GPA in case of guest page fault
    );

    //# Context Directory Walker
    rv_iommu_cdw_ext #(
        .axi_req_t          (axi_req_t ),
        .axi_rsp_t          (axi_rsp_t )
    ) i_rv_iommu_cdw_ext (
        .clk_i                  (clk_i              ),  // Clock
        .rst_ni                 (rst_ni             ),  // Asynchronous reset active low
        
        // Error signaling
        .cdw_active_o           (cdw_active         ),  // Set when CDW is walking memory
        .cdw_error_o            (cdw_error          ),  // set when an error occurred
        .cause_code_o           (cdw_cause_code     ),  // Fault code as defined by IOMMU and Priv Spec

        // DC config checks
        .caps_ats_i             (capabilities_i.ats.q       ),
        .caps_t2gpa_i           (capabilities_i.t2gpa.q     ),
        .caps_pd20_i            (capabilities_i.pd20.q      ),
        .caps_pd17_i            (capabilities_i.pd17.q      ),
        .caps_pd8_i             (capabilities_i.pd8.q       ),
        .caps_sv32_i            (capabilities_i.sv32.q      ),
        .caps_sv39_i            (capabilities_i.sv39.q      ),
        .caps_sv48_i            (capabilities_i.sv48.q      ), 
        .caps_sv57_i            (capabilities_i.sv57.q      ),
        .fctl_gxl_i             (fctl_i.gxl.q               ),
        .caps_sv32x4_i          (capabilities_i.sv32x4.q    ),
        .caps_sv39x4_i          (capabilities_i.sv39x4.q    ),
        .caps_sv48x4_i          (capabilities_i.sv48x4.q    ),
        .caps_sv57x4_i          (capabilities_i.sv57x4.q    ),
        .caps_msi_flat_i        (capabilities_i.msi_flat.q  ),
        .caps_amo_hwad_i        (capabilities_i.amo_hwad.q  ),
        .caps_end_i             (capabilities_i.endi.q      ),
        .fctl_be_i              (fctl_i.be.q                ),

        // CDW memory interface
        .mem_resp_i             (cdw_axi_resp_i ),      // Response port from memory
        .mem_req_o              (cdw_axi_req_o  ),      // Request port to memory

        // Update logic
        .update_dc_o            (ddtc_update    ),
        .up_did_o               (ddtc_up_did    ),
        .up_dc_content_o        (ddtc_up_content),

        // CDCs tags
        .req_did_i              (did_i          ),      // device ID associated with request

        // from DDTC, to monitor misses
        .ddtc_access_i          (ddtc_access    ),
        .ddtc_hit_i             (ddtc_lu_hit    ),

        // from regmap
        .ddtp_ppn_i             (ddtp_i.ppn.q       ),  // PPN from ddtp register
        .ddtp_mode_i            (ddtp_i.iommu_mode.q)   // DDT levels and IOMMU mode
    );

    //# Translation logic
    always_comb begin : translation

        ddtc_access         = 1'b0;
        en_1S               = 1'b0;
        en_2S               = 1'b0;
        gscid               = '0;
        pscid               = '0;
        iosatp_ppn          = '0;
        iohgatp_ppn         = '0;
        iotlb_access        = 1'b0;
        cause_code          = '0;
        trans_error         = 1'b0;
        is_msi_o            = 1'b0;
        trans_valid_o       = 1'b0;
        spaddr_o   = '0;
        report_always       = 1'b0;

        // A translation is triggered by setting req_trans_i
        if (req_trans_i) begin
    
            //# Input Checks
            // "If ddtp.iommu_mode == Off then stop and report "All inbound transactions disallowed" (cause = 256)."
            if (ddtp_i.iommu_mode.q == 4'b0000) begin
                cause_code    = rv_iommu::ALL_INB_TRANSACTIONS_DISALLOWED;
                trans_error   = 1'b1;
                report_always   = 1'b1;
            end

            // "If ddtp.iommu_mode == Bare and any of the following conditions (*) hold then stop and report "Transaction type disallowed" (cause = 260)."
            else if (ddtp_i.iommu_mode.q == 4'b0001) begin
                
                // "(*) If the transaction is a translated request or a PCIe ATS request"
                if (is_translated || is_pcie_tr_req) begin
                    cause_code    = rv_iommu::TRANS_TYPE_DISALLOWED;
                    trans_error   = 1'b1;
                    report_always   = 1'b1;
                end

                // " else the translation process is completed with the IOVA as the translated address"
                else begin
                    trans_valid_o       = 1'b1;
                    spaddr_o   = iova_i[riscv::PLEN-1:0];
                end
            end

            // This implementation will support MSI address translation, so DC always is presented in extended format

            // "If the device_id is wider than supported by the IOMMU, then stop and report "Transaction type disallowed" (cause = 260)."
            else if ((ddtp_i.iommu_mode.q == 4'b0011 && (|did_i[23:15])) || (ddtp_i.iommu_mode.q == 4'b0010 && (|did_i[23:6]))) begin
                cause_code = rv_iommu::TRANS_TYPE_DISALLOWED;
                trans_error   = 1'b1;
                report_always   = 1'b1;
            end

            // IOMMU is not in bare mode and no errors ocurred. Lookup DDTC
            else ddtc_access = 1'b1;
        end

        //# DDTC Lookup
        // Access to DDTC and PDTC is automatically triggered when setting req_trans_i if no fault is generated
        // If hit flag is set in the same cycle, we have a DDTC instantaneous hit
        if (ddtc_lu_hit) begin

            // "If any of the following conditions hold then stop and report "Transaction type disallowed" (cause = 260)."
            if (((is_translated || is_pcie_tr_req) && !ddtc_lu_content.tc.en_ats)) begin

                cause_code  = rv_iommu::TRANS_TYPE_DISALLOWED;
                trans_error = 1'b1;
            end

            // avoid triggering a CDW walk for a PC or a PTW walk when the previous fault occurs 
            else begin

                // Translated request
                if (is_translated) begin

                    // When DC.tc.T2GPA = 0, translated requests are performed using an SPA. Translation process is complete
                    if (!ddtc_lu_content.tc.t2gpa) begin
                        trans_valid_o       = 1'b1;
                        spaddr_o   = iova_i[riscv::PLEN-1:0];
                    end

                    // If DC.tc.T2GPA = 1, translated requests are performed using a GPA. The IOMMU performs second-stage translation
                    else begin
                        // Stage 1 Bare
                        en_2S           = ~second_stage_is_bare;
                        gscid           = ddtc_lu_content.iohgatp.gscid;
                        // PSCID not used since Stage 1 is Bare
                        iohgatp_ppn     = ddtc_lu_content.iohgatp.ppn;
                        // iosatp not used since Stage 1 is Bare
                        iotlb_access    = 1'b1;
                    end
                end

                // Untranslated request
                else begin
                    
                    // No Process Context
                    if (!ddtc_lu_content.tc.pdtv) begin
                        en_1S           = ~first_stage_is_bare;
                        en_2S           = ~second_stage_is_bare;
                        gscid           = ddtc_lu_content.iohgatp.gscid;
                        pscid           = ddtc_lu_content.ta.pscid;
                        iohgatp_ppn     = ddtc_lu_content.iohgatp.ppn;
                        iosatp_ppn      = ddtc_lu_content.fsc.ppn;
                        iotlb_access    = 1'b1;
                    end

                    // Process Context associated
                    // Raise fault since this module does not support PCs
                    else begin
                        cause_code  = rv_iommu::TRANS_TYPE_DISALLOWED;
                        trans_error = 1'b1;
                    end
                end
            end

            //# IOTLB Lookup
            if (iotlb_lu_hit) begin
                
                trans_valid_o       = 1'b1;

                //# MSI addr entry
                if (iotlb_lu_is_msi && msi_enabled) begin
                    is_msi_o            = 1'b1;
                    // MSI PTEs contain the PPN in the same position as normal PTEs
                    spaddr_o   = {iotlb_lu_2S_content.ppn, iova_i[11:0]};
                end

                //# Normal entry
                // INFO: IOTLB should not have entries with both stages disabled and MSI flag clear. However, we double-check
                else if (en_1S || en_2S) begin
                    /*
                    A fault is generated if:
                        - A bit is not set (checked in PTW);
                        - Page is not readable (checked in PTW);
                        - (1): Transaction is a store and page has not write permissions (D bit checked in PTW);
                        - (2): Transaction is read-for-execute and page has not X permissions;
                        - (3): U-mode transaction and PTE has U=0;
                    */
                    if  ((is_store && (!iotlb_lu_1S_content.w && en_1S)                                     ) ||        // (1)
                         (is_rx && (!iotlb_lu_1S_content.x && en_1S)                                        ) ||        // (2)
                         (!iotlb_lu_1S_content.u && en_1S                                                   )           // (3)
                        ) begin
                            if (is_store)   cause_code = rv_iommu::STORE_PAGE_FAULT;
                            else            cause_code = rv_iommu::LOAD_PAGE_FAULT;
                            trans_error     = 1'b1;
                            trans_valid_o   = 1'b0;
                    end

                    else if ((is_store && (!iotlb_lu_2S_content.w && en_2S)  ) ||    // (1)
                             (is_rx && (!iotlb_lu_2S_content.x && en_2S)     )       // (2)
                            ) begin
                            if (is_store)   cause_code = rv_iommu::STORE_GUEST_PAGE_FAULT;
                            else            cause_code = rv_iommu::LOAD_GUEST_PAGE_FAULT;
                            trans_error     = 1'b1;
                            trans_valid_o   = 1'b0;
                    end 

                    //# Address Translation Found
                    else begin
                        
                        spaddr_o = {((en_2S) ? iotlb_lu_2S_content.ppn : iotlb_lu_1S_content.ppn), iova_i[11:0]};

                        // Apply superpage cases
                        if (en_1S && en_2S) begin
                            case ({iotlb_lu_1S_2M, iotlb_lu_1S_1G, iotlb_lu_2S_2M, iotlb_lu_2S_1G})

                                // 1-S: 4k | 2-S: 2M:   {PPN[2], PPN[1],  GPPN[0], OFF}
                                4'b0010:    spaddr_o[20:12] = iotlb_lu_1S_content.ppn[20:12];

                                // 1-S: 2M | 2-S: 2M:   {PPN[2], PPN[1],  VPN[0],  OFF}
                                // 1-S: 1G | 2-S: 2M:   {PPN[2], PPN[1],  VPN[0],  OFF}
                                4'b1010, 4'b0110:   spaddr_o[20:12] = iova_i[20:12];

                                // 1-S: 4k | 2-S: 1G:   {PPN[2], GPPN[1], GPPN[0], OFF}
                                4'b0001:    spaddr_o[29:12] = iotlb_lu_1S_content.ppn[29:12];

                                // 1-S: 1G | 2-S: 1G:   {PPN[2], VPN[1],  VPN[0],  OFF}
                                4'b0101:    spaddr_o[29:12] = iova_i[29:12];

                                // 1-S: 2M | 2-S: 1G:   {PPN[2], GPPN[1], VPN[0],  OFF}
                                4'b1001:    spaddr_o[29:12] = {iotlb_lu_1S_content.ppn[29:21], iova_i[20:12]};
                                
                                default:;
                                    // 1-S: 4k | 2-S: 4k:   {PPN[2], PPN[1],  PPN[0],  OFF}
                                    // 1-S: 2M | 2-S: 4k:   {PPN[2], PPN[1],  PPN[0],  OFF}
                                    // 1-S: 1G | 2-S: 4k:   {PPN[2], PPN[1],  PPN[0],  OFF}
                            endcase
                        end

                        else begin
                            if (iotlb_lu_2S_1G || iotlb_lu_1S_1G)   spaddr_o[29:12] = iova_i[29:12];
                            if (iotlb_lu_2S_2M || iotlb_lu_1S_2M)   spaddr_o[20:12] = iova_i[20:12];
                        end
                    end
                end

                /*
                    # Note about IOPMP faults for translated IOVAs:
                    IOPMP access faults are reported as failing AXI transactions. After translating the IOVA,
                    the AXI transaction continues without IOMMU intervention (data is opaque to the IOMMU).
                    If the translated physical address violates an IOPMP check, the requesting device will be
                    responded by the IOPMP with an AXI error.
                */
            end

            // No stage is enabled and input address does not correspond to a MSI address
            // (This condition and an IOTLB hit should be mutually exclusive)
            // Input address is bypassed
            if (is_bare_translation) begin
                trans_valid_o     = 1'b1;
                spaddr_o = iova_i[riscv::PLEN-1:0];
            end
        end

        //# Check for errors
        // If we had to walk memory is because we had a miss. As we had an exception,
        // the corresponding cache/TLB was not updated, and translation was never set to valid
        if (ptw_error || cdw_error || msi_write_error_i) begin
            cause_code    = (cdw_error) ? cdw_cause_code : ptw_cause_code;
            trans_error   = 1'b1;
        end
    end

endmodule